//-- sv_mi_common_pkg.sv: Package for common mi fifo verification
//-- Copyright (C) 2021 CESNET z. s. p. o.
//-- Author(s): Tomáš Beneš <xbenes55@stud.fit.vutbr.cz>
//--
//-- SPDX-License-Identifier: BSD-3-Clause 

package sv_mi_common_pkg; 

    `include "mi_common_scoreboard.sv"

endpackage
