/*
 * file       : pkg.sv
 * Copyright (C) 2021 CESNET z. s. p. o.
 * description: RESET packages 
 * date       : 2021
 * author     : Radek Iša <isa@cesnet.cz>
 *
 * SPDX-License-Identifier: BSD-3-Clause
*/


`ifndef RESET_PKG
`define RESET_PKG

package reset;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "sync.sv"
    `include "config.sv"

    `include "sequence_item.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent.sv"
    `include "sequence.sv"

    //enviroment with more resets
    `include "env_driver.sv"
    `include "low_sequence.sv"
    `include "env_config.sv"
    `include "env.sv"
endpackage


`endif
