//-- pkg.sv
//-- Copyright (C) 2022 CESNET z. s. p. o.
//-- Author(s): Daniel Kriz <danielkriz@cesnet.cz>

//-- SPDX-License-Identifier: BSD-3-Clause


`ifndef INFO_PKG
`define INFO_PKG

package uvm_dma_ll_info;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "watchdog.sv"

endpackage

`endif
