//-- pkg.sv: Package for AXI interface
//-- Copyright (C) 2022 CESNET z. s. p. o.
//-- Author(s): Daniel Kříž <xkrizd01@vutbr.cz>

//-- SPDX-License-Identifier: BSD-3-Clause 

`ifndef AXI_PKG
`define AXI_PKG

package uvm_axi;
    
    `include "uvm_macros.svh"
    import uvm_pkg::*;
   
    `include "config.sv"
    `include "sequence_item.sv"
    `include "sequencer.sv"
    `include "sequence.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent.sv"
endpackage

`endif
