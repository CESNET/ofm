/*!
 * \file sv_fifox_cov_pkg.sv
 * \brief Coverages package for verification
 * \author Tomáš Beneš <xbenes55@stud.fit.vutbr.cz>
 * \date 2016
*/
/*
 * SPDX-License-Identifier: BSD-3-Clause
*/

package sv_fifox_cov_pkg;
  `include "fifox_in_cov.sv"
  `include "fifox_out_cov.sv"
endpackage
