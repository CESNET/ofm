/*!
 * \file scoreboard.sv
 * \brief Score Board
 * \author Lukas Kekely <kekely@cesnet.cz>
 * \date 2016
 */
 /*
 * Copyright (C) 2015 CESNET
 *
 * LICENSE TERMS
 *
 * SPDX-License-Identifier: BSD-3-Clause
 *
 */

import sv_common_pkg::*;
import sv_flu_pkg::*;



class ScoreboardDriverCbs extends DriverCbs;

    TransactionTable #(0) sc_table;


    function new (TransactionTable #(0) sc_table);
        this.sc_table = sc_table;
    endfunction

    virtual task post_tx(Transaction transaction, string inst);
        sc_table.add(transaction);
    endtask

endclass : ScoreboardDriverCbs



class ScoreboardMonitorCbs extends MonitorCbs;

    TransactionTable #(0) sc_table;


    function new (TransactionTable #(0) sc_table);
        this.sc_table = sc_table;
    endfunction

    virtual task post_rx(Transaction transaction, string inst);
        bit status=0;
        sc_table.remove(transaction, status);
        if (status==0)begin
            $write("Unknown transaction received from monitor %d\n", inst);
            $timeformat(-9, 3, " ns", 8);
            $write("Time: %t\n", $time);
            transaction.display();
            sc_table.display();
            $stop;
        end;
    endtask

endclass : ScoreboardMonitorCbs



class Scoreboard;

    TransactionTable #(0) scoreTable;
    ScoreboardMonitorCbs  monitorCbs;
    ScoreboardDriverCbs   driverCbs;


    function new ();
        this.scoreTable = new;
        this.monitorCbs = new(scoreTable);
        this.driverCbs  = new(scoreTable);
    endfunction

    task display();
        scoreTable.display();
    endtask
  
endclass : Scoreboard
