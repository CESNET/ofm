//-- pkg.sv: Package for environment
//-- Copyright (C) 2022 CESNET z. s. p. o.
//-- Author:   Daniel Kříž <xkrizd01@vutbr.cz>

//-- SPDX-License-Identifier: BSD-3-Clause

`ifndef FIFOX_ENV_SV
`define FIFOX_ENV_SV

package uvm_pipe;
    
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "scoreboard.sv"
    `include "env.sv"
    `include "model.sv"

endpackage

`endif
