/*
 * pkg.sv scoremoard package 
 * Copyright (C) 2020 CESNET z. s. p. o.
 * Author(s): Radek Iša <isa@cesnet.cz>
 * SPDX-License-Identifier: BSD-3-Clause
 */

package scoreboard;
    `include "data.sv"
    `include "cbs.sv"
    `include "sc.sv"
endpackage
