-- buffer.vhd:
-- Copyright (C) 2019 CESNET z. s. p. o.
-- Author(s): Jakub Cabal <cabal@cesnet.cz>
--
-- SPDX-License-Identifier: BSD-3-Clause

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.math_pack.all;
use work.type_pack.all;

entity RX_MAC_LITE_BUFFER is
    generic(
        REGIONS        : natural := 4;
        REGION_SIZE    : natural := 8;
        BLOCK_SIZE     : natural := 8;
        ITEM_WIDTH     : natural := 8;
        META_WIDTH     : natural := 16;
        META_ALIGN2SOF : boolean := True;
        DFIFO_ITEMS    : natural := 512;
        MFIFO_ITEMS    : natural := 32;
        MFIFO_RAM_TYPE : string  := "LUT";
        DEVICE         : string  := "STRATIX10"
    );
   port(
        -- =====================================================================
        -- INPUT INTERFACES
        -- =====================================================================
        -- CLOCK AND RESET
        -- ---------------------------------------------------------------------
        RX_CLK          : in  std_logic;
        RX_RESET        : in  std_logic;

        -- MFB BUS WITH METADATA AND ERROR FLAG (ALIGNED TO EOF)
        -- ---------------------------------------------------------------------
        RX_DATA         : in  std_logic_vector(REGIONS*REGION_SIZE*BLOCK_SIZE*ITEM_WIDTH-1 downto 0);
        RX_SOF_POS      : in  std_logic_vector(REGIONS*max(1,log2(REGION_SIZE))-1 downto 0);
        RX_EOF_POS      : in  std_logic_vector(REGIONS*max(1,log2(REGION_SIZE*BLOCK_SIZE))-1 downto 0);
        RX_SOF          : in  std_logic_vector(REGIONS-1 downto 0);
        RX_EOF          : in  std_logic_vector(REGIONS-1 downto 0);
        RX_ERROR        : in  std_logic_vector(REGIONS-1 downto 0);
        RX_METADATA     : in  slv_array_t(REGIONS-1 downto 0)(META_WIDTH-1 downto 0);
        RX_SRC_RDY      : in  std_logic;

        -- STATISTICS OUTPUT
        -- ---------------------------------------------------------------------
        BUFFER_STATUS   : out std_logic_vector(2-1 downto 0);
        STAT_BUFFER_OVF : out std_logic_vector(REGIONS-1 downto 0);
        STAT_DISCARD    : out std_logic_vector(REGIONS-1 downto 0);
        STAT_METADATA   : out slv_array_t(REGIONS-1 downto 0)(META_WIDTH-1 downto 0);
        STAT_VALID      : out std_logic_vector(REGIONS-1 downto 0);

        -- =====================================================================
        -- OUTPUT INTERFACES
        -- =====================================================================
        -- CLOCK AND RESET
        -- ---------------------------------------------------------------------
        TX_CLK          : in  std_logic;
        TX_RESET        : in  std_logic;

        -- MFB BUS
        -- ---------------------------------------------------------------------
        TX_MFB_DATA     : out std_logic_vector(REGIONS*REGION_SIZE*BLOCK_SIZE*ITEM_WIDTH-1 downto 0);
        TX_MFB_SOF_POS  : out std_logic_vector(REGIONS*max(1,log2(REGION_SIZE))-1 downto 0);
        TX_MFB_EOF_POS  : out std_logic_vector(REGIONS*max(1,log2(REGION_SIZE*BLOCK_SIZE))-1 downto 0);
        TX_MFB_SOF      : out std_logic_vector(REGIONS-1 downto 0);
        TX_MFB_EOF      : out std_logic_vector(REGIONS-1 downto 0);
        TX_MFB_SRC_RDY  : out std_logic;
        TX_MFB_DST_RDY  : in  std_logic;

        -- MVB BUS
        -- ---------------------------------------------------------------------
        TX_MVB_DATA     : out std_logic_vector(REGIONS*META_WIDTH-1 downto 0);
        TX_MVB_VLD      : out std_logic_vector(REGIONS-1 downto 0);
        TX_MVB_SRC_RDY  : out std_logic;
        TX_MVB_DST_RDY  : in  std_logic
    );
end entity;

architecture FULL of RX_MAC_LITE_BUFFER is

    constant SOF_INDEX_WIDTH : natural := log2(REGIONS);
    constant MBUF_WIDTH      : natural := META_WIDTH+SOF_INDEX_WIDTH+1+1;

    type fsm_t is (st_idle, st_recovery);

    signal s_inc_frame          : std_logic_vector(REGIONS downto 0);
    signal s_inc_frame_reg      : std_logic;
    signal s_whole_frame        : std_logic_vector(REGIONS-1 downto 0);

    signal fsm_pst              : fsm_t;
    signal fsm_nst              : fsm_t;
    signal s_wait_for_recovery  : std_logic;
    signal s_rx_eof_removed     : std_logic_vector(REGIONS-1 downto 0);
    signal s_rx_src_rdy_clear   : std_logic;
    signal s_rx_recovered       : std_logic;

    signal s_rx_data_reg        : std_logic_vector(REGIONS*REGION_SIZE*BLOCK_SIZE*ITEM_WIDTH-1 downto 0);
    signal s_rx_sof_pos_reg     : std_logic_vector(REGIONS*max(1,log2(REGION_SIZE))-1 downto 0);
    signal s_rx_eof_pos_reg     : std_logic_vector(REGIONS*max(1,log2(REGION_SIZE*BLOCK_SIZE))-1 downto 0);
    signal s_rx_sof_reg         : std_logic_vector(REGIONS-1 downto 0);
    signal s_rx_eof_reg         : std_logic_vector(REGIONS-1 downto 0);
    signal s_rx_error_reg       : std_logic_vector(REGIONS-1 downto 0);
    signal s_rx_metadata_reg    : slv_array_t(REGIONS-1 downto 0)(META_WIDTH-1 downto 0);
    signal s_rx_src_rdy_reg     : std_logic;
    signal s_rx_eof_removed_reg : std_logic_vector(REGIONS-1 downto 0);
    signal s_rx_recovered_reg   : std_logic;
    signal s_whole_frame_reg    : std_logic_vector(REGIONS-1 downto 0);

    signal s_rx_stop_reg        : std_logic;
    signal s_rx_stop_reg2       : std_logic;

    signal s_full_flag          : std_logic;
    signal s_stop_reg           : std_logic;
    signal s_stop_flag          : std_logic;

    signal s_dbuf_wr            : std_logic;
    signal s_dbuf_rdy           : std_logic;
    signal s_dbuf_full          : std_logic;
    signal s_dbuf_discard       : std_logic_vector(REGIONS-1 downto 0);
    signal s_dbuf_force_discard : std_logic;

    signal s_last_sof           : std_logic_vector(REGIONS-1 downto 0);
    signal s_dist_sof_index     : slv_array_t(REGIONS downto 0)(SOF_INDEX_WIDTH-1 downto 0);
    signal s_dist_sof_liw       : std_logic_vector(REGIONS downto 0);
    signal s_dist_sof_index_fix : slv_array_t(REGIONS-1 downto 0)(SOF_INDEX_WIDTH-1 downto 0);
    signal s_dist_sof_liw_fix   : std_logic_vector(REGIONS-1 downto 0);
    signal s_fake_item          : std_logic_vector(REGIONS-1 downto 0);
    signal s_fake_item_vld      : std_logic_vector(REGIONS-1 downto 0);
    signal s_fake_item_src_rdy  : std_logic;

    signal s_meta_vld           : std_logic_vector(REGIONS-1 downto 0);
    signal s_meta_src_rdy       : std_logic;

    signal s_mbuf_din           : slv_array_t(REGIONS-1 downto 0)(MBUF_WIDTH-1 downto 0);
    signal s_mbuf_vld           : std_logic_vector(REGIONS-1 downto 0);
    signal s_mbuf_src_rdy       : std_logic;
    signal s_mbuf_status        : std_logic_vector(log2(MFIFO_ITEMS) downto 0);
    signal s_mbuf_afull         : std_logic;
    signal s_mbuf_afull_reg     : std_logic;
    signal s_mbuf_afull_reg2    : std_logic;
    signal s_mbuf_dout_ser      : std_logic_vector(REGIONS*MBUF_WIDTH-1 downto 0);
    signal s_mbuf_dout          : slv_array_t(REGIONS-1 downto 0)(MBUF_WIDTH-1 downto 0);
    signal s_mbuf_mvb_data      : slv_array_t(REGIONS-1 downto 0)(META_WIDTH-1 downto 0);
    signal s_mbuf_mvb_new_pos   : slv_array_t(REGIONS-1 downto 0)(SOF_INDEX_WIDTH-1 downto 0);
    signal s_mbuf_mvb_new_liw   : std_logic_vector(REGIONS-1 downto 0);
    signal s_mbuf_mvb_fake      : std_logic_vector(REGIONS-1 downto 0);
    signal s_mbuf_mvb_vld       : std_logic_vector(REGIONS-1 downto 0);
    signal s_mbuf_mvb_src_rdy   : std_logic;
    signal s_mbuf_mvb_dst_rdy   : std_logic;
  
begin

    -- -------------------------------------------------------------------------
    --  FRAME STATE LOGIC
    -- -------------------------------------------------------------------------

    inc_frame_g : for r in 0 to REGIONS-1 generate
        s_inc_frame(r+1) <= (RX_SOF(r) and not RX_EOF(r) and not s_inc_frame(r)) or
                            (RX_SOF(r) and RX_EOF(r) and s_inc_frame(r)) or
                            (not RX_SOF(r) and not RX_EOF(r) and s_inc_frame(r));
    end generate;

    inc_frame_last_reg_p : process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            if (RX_RESET = '1') then
                s_inc_frame(0)  <= '0';
                s_inc_frame_reg <= '0';
            elsif (RX_SRC_RDY = '1') then
                s_inc_frame(0)  <= s_inc_frame(REGIONS);
                s_inc_frame_reg <= s_inc_frame(REGIONS); -- register duplication for better timing
            end if;
        end if;
    end process;

    s_whole_frame <= RX_SOF and RX_EOF and not s_inc_frame(REGIONS-1 downto 0);

    -- -------------------------------------------------------------------------
    --  AFTER BUFFER OVERFULL RECOVERY LOGIC
    -- -------------------------------------------------------------------------

    process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            fsm_pst <= fsm_nst;
            if (RX_RESET = '1') then
                fsm_pst <= st_idle;
            end if;
        end if;
    end process;

    process (all)
    begin
        fsm_nst <= fsm_pst;
        case (fsm_pst) is
            when st_idle =>
                s_wait_for_recovery <= '0';
                if (s_rx_stop_reg = '0' and s_rx_stop_reg2 = '1') then
                    fsm_nst <= st_recovery;
                end if;

            when st_recovery =>
                s_wait_for_recovery <= '1';
                if (s_rx_recovered = '1') then
                    fsm_nst <= st_idle;
                end if;
        end case;
    end process;

    process (all)
    begin
        s_rx_eof_removed <= (others => '0');
        for r in 0 to REGIONS-1 loop
            if (RX_EOF(r) = '1') then
                s_rx_eof_removed(r) <= RX_SRC_RDY and s_wait_for_recovery and s_inc_frame_reg;
                exit;
            end if;
        end loop;
    end process;

    s_rx_src_rdy_clear <= not (or RX_SOF) and s_inc_frame_reg and s_wait_for_recovery;
    s_rx_recovered <= ((RX_SRC_RDY and (or RX_EOF)) or (not RX_SRC_RDY and not s_inc_frame_reg)) and s_wait_for_recovery;

    -- -------------------------------------------------------------------------
    --  REGISTER STAGE
    -- -------------------------------------------------------------------------

    process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            s_rx_data_reg        <= RX_DATA;
            s_rx_sof_pos_reg     <= RX_SOF_POS;
            s_rx_eof_pos_reg     <= RX_EOF_POS;
            s_rx_sof_reg         <= RX_SOF;
            s_rx_eof_reg         <= RX_EOF and not s_rx_eof_removed;
            s_rx_error_reg       <= RX_ERROR;
            s_rx_metadata_reg    <= RX_METADATA;
            s_rx_eof_removed_reg <= s_rx_eof_removed;
            s_whole_frame_reg    <= s_whole_frame;
        end if;
    end process;
    
    process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            if (RX_RESET = '1') then
                s_rx_src_rdy_reg   <= '0';
                s_rx_recovered_reg <= '0';
            else
                s_rx_src_rdy_reg   <= RX_SRC_RDY and not s_rx_src_rdy_clear;
                s_rx_recovered_reg <= s_rx_recovered;
            end if;
        end if;
    end process;

    process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            if (RX_RESET = '1') then
                s_rx_stop_reg  <= '0';
                s_rx_stop_reg2 <= '0';
            else
                s_rx_stop_reg  <= s_full_flag;
                s_rx_stop_reg2 <= s_rx_stop_reg;
            end if;
        end if;
    end process;

    -- -------------------------------------------------------------------------
    --  FIFOs CONTROL LOGIC
    -- -------------------------------------------------------------------------

    s_full_flag <= s_dbuf_full or s_mbuf_afull_reg2;

    stop_reg_p : process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            if (RX_RESET = '1') then
                s_stop_reg <= '0';
            elsif (s_full_flag = '1') then
                s_stop_reg <= '1';
            elsif (s_rx_recovered_reg = '1') then
                s_stop_reg <= '0';  
            end if;
        end if;
    end process;

    s_stop_flag <= s_full_flag or (s_stop_reg and not s_rx_recovered_reg);

    s_dbuf_wr            <= s_rx_src_rdy_reg;
    s_dbuf_full          <= not s_dbuf_rdy;
    s_dbuf_discard       <= s_rx_error_reg;
    s_dbuf_force_discard <= s_stop_flag;

    buffer_status_reg_p : process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            BUFFER_STATUS(0) <= s_mbuf_afull_reg2 and s_rx_src_rdy_reg;
            BUFFER_STATUS(1) <= s_dbuf_full and s_rx_src_rdy_reg;
        end if;
    end process;

    -- -------------------------------------------------------------------------
    --  STATISTICS OUTPUT
    -- -------------------------------------------------------------------------

    process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            STAT_BUFFER_OVF <= (s_rx_src_rdy_reg and s_rx_eof_reg and s_stop_flag) or s_rx_eof_removed_reg;
            STAT_DISCARD    <= (s_rx_src_rdy_reg and s_rx_eof_reg and (s_rx_error_reg or s_stop_flag)) or s_rx_eof_removed_reg;
            STAT_METADATA   <= s_rx_metadata_reg;
            STAT_VALID      <= (s_rx_src_rdy_reg and s_rx_eof_reg) or s_rx_eof_removed_reg;
            if (RX_RESET = '1') then
                STAT_VALID <= (others => '0');
            end if;
        end if;
    end process;

    -- -------------------------------------------------------------------------
    --  DATA and META BUFFER
    -- -------------------------------------------------------------------------

    dbuf_i : entity work.MFB_PD_ASFIFO
    generic map(
        REGIONS     => REGIONS,
        REGION_SIZE => REGION_SIZE,
        BLOCK_SIZE  => BLOCK_SIZE,
        ITEM_WIDTH  => ITEM_WIDTH,
        ITEMS       => DFIFO_ITEMS,
        DEVICE      => DEVICE
    )
    port map(
        RX_CLK           => RX_CLK,
        RX_RESET         => RX_RESET,

        RX_DATA          => s_rx_data_reg,
        RX_SOF_POS       => s_rx_sof_pos_reg,
        RX_EOF_POS       => s_rx_eof_pos_reg,
        RX_SOF           => s_rx_sof_reg,
        RX_EOF           => s_rx_eof_reg,
        RX_SRC_RDY       => s_dbuf_wr,
        RX_DST_RDY       => s_dbuf_rdy,

        RX_DISCARD       => s_dbuf_discard,
        RX_FORCE_DISCARD => s_dbuf_force_discard,
        STATUS           => open,

        TX_CLK           => TX_CLK,
        TX_RESET         => TX_RESET,
        
        TX_DATA          => TX_MFB_DATA,
        TX_SOF_POS       => TX_MFB_SOF_POS,
        TX_EOF_POS       => TX_MFB_EOF_POS,
        TX_SOF           => TX_MFB_SOF,
        TX_EOF           => TX_MFB_EOF,
        TX_SRC_RDY       => TX_MFB_SRC_RDY,
        TX_DST_RDY       => TX_MFB_DST_RDY
    );

    dist_sof_g: if META_ALIGN2SOF generate
        last_sof_p : process (all)
        begin
            s_last_sof <= (others => '0');
            for i in REGIONS-1 downto 0 loop
                if (s_rx_sof_reg(i) = '1') then
                    s_last_sof(i) <= '1';
                    exit;
                end if;
            end loop;
        end process;

        dist_sof_g : for i in 0 to REGIONS-1 generate
            dist_sof_p : process (all)
            begin
                if (s_rx_sof_reg(i) = '1') then
                    s_dist_sof_index(i+1) <= std_logic_vector(to_unsigned(i,SOF_INDEX_WIDTH));
                    s_dist_sof_liw(i+1)   <= s_last_sof(i);
                else
                    s_dist_sof_index(i+1) <= s_dist_sof_index(i);
                    s_dist_sof_liw(i+1)   <= s_dist_sof_liw(i);
                end if;
            end process;
        end generate;

        dist_sof_fix_g : for i in 0 to REGIONS-1 generate
            dist_sof_fix_p : process (all)
            begin
                if (s_whole_frame_reg(i) = '1') then
                    s_dist_sof_index_fix(i) <= std_logic_vector(to_unsigned(i,SOF_INDEX_WIDTH));
                    s_dist_sof_liw_fix(i)   <= s_last_sof(i);
                else
                    s_dist_sof_index_fix(i) <= s_dist_sof_index(i);
                    s_dist_sof_liw_fix(i)   <= s_dist_sof_liw(i);
                end if;
            end process;
        end generate;

        dist_sof_reg_p : process (RX_CLK)
        begin
            if (rising_edge(RX_CLK)) then
                if (s_rx_src_rdy_reg = '1') then
                    s_dist_sof_index(0) <= s_dist_sof_index(REGIONS);
                    s_dist_sof_liw(0)   <= s_dist_sof_liw(REGIONS);
                end if;
            end if;
        end process;

        s_fake_item         <= s_rx_error_reg or s_stop_flag;
        s_fake_item_vld     <= s_dist_sof_liw_fix and s_rx_eof_reg and s_rx_src_rdy_reg;
        s_fake_item_src_rdy <= or s_fake_item_vld;
    else generate
        s_dist_sof_index_fix <= (others => (others => '0'));
        s_dist_sof_liw_fix   <= (others => '0');

        s_fake_item         <= (others => '0');
        s_fake_item_vld     <= (others => '0');
        s_fake_item_src_rdy <= '0';
    end generate;

    s_meta_vld <= s_rx_eof_reg and not s_rx_error_reg and not s_stop_flag and s_rx_src_rdy_reg;
    s_meta_src_rdy <= or s_meta_vld;

    mbuf_din_g : for i in 0 to REGIONS-1 generate
        s_mbuf_din(i) <= s_rx_metadata_reg(i) & s_dist_sof_index_fix(i) & s_dist_sof_liw_fix(i) & s_fake_item(i);
    end generate;

    s_mbuf_vld     <= s_meta_vld or s_fake_item_vld;
    s_mbuf_src_rdy <= s_meta_src_rdy or s_fake_item_src_rdy;

    mbuf_i : entity work.MVB_ASFIFOX
    generic map(
        MVB_ITEMS      => REGIONS,
        MVB_ITEM_WIDTH => MBUF_WIDTH,
        FIFO_ITEMS     => MFIFO_ITEMS,
        RAM_TYPE       => MFIFO_RAM_TYPE,
        FWFT_MODE      => True,
        OUTPUT_REG     => True,
        DEVICE         => DEVICE
    )
    port map(
        RX_CLK     => RX_CLK,
        RX_RESET   => RX_RESET,
        RX_DATA    => slv_array_ser(s_mbuf_din,REGIONS,MBUF_WIDTH),
        RX_VLD     => s_mbuf_vld,
        RX_SRC_RDY => s_mbuf_src_rdy,
        RX_DST_RDY => open,
        RX_AFULL   => open,
        RX_STATUS  => s_mbuf_status,

        TX_CLK     => TX_CLK,
        TX_RESET   => TX_RESET,
        TX_DATA    => s_mbuf_dout_ser,
        TX_VLD     => s_mbuf_mvb_vld,
        TX_SRC_RDY => s_mbuf_mvb_src_rdy,
        TX_DST_RDY => s_mbuf_mvb_dst_rdy
    );

    process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            if (RX_RESET = '1') then
                s_mbuf_afull <= '1';
            elsif (unsigned(s_mbuf_status) >= (MFIFO_ITEMS-6)) then
                s_mbuf_afull <= '1';
            elsif (unsigned(s_mbuf_status) < (MFIFO_ITEMS-MFIFO_ITEMS/4)) then
                s_mbuf_afull <= '0';
            end if;
        end if;
    end process;

    mbuf_afull_reg_p : process (RX_CLK)
    begin
        if (rising_edge(RX_CLK)) then
            if (RX_RESET = '1') then
                s_mbuf_afull_reg  <= '1';
                s_mbuf_afull_reg2 <= '1';
            else
                s_mbuf_afull_reg  <= s_mbuf_afull;
                s_mbuf_afull_reg2 <= s_mbuf_afull_reg;
            end if;
        end if;
    end process;

    s_mbuf_dout <= slv_array_downto_deser(s_mbuf_dout_ser,REGIONS,MBUF_WIDTH);

    mbuf_mvb_g : for i in 0 to REGIONS-1 generate
        s_mbuf_mvb_data(i)    <= s_mbuf_dout(i)(MBUF_WIDTH-1 downto 2+SOF_INDEX_WIDTH);
        s_mbuf_mvb_new_pos(i) <= s_mbuf_dout(i)(2+SOF_INDEX_WIDTH-1 downto 2);
        s_mbuf_mvb_new_liw(i) <= s_mbuf_dout(i)(1);
        s_mbuf_mvb_fake(i)    <= s_mbuf_dout(i)(0);
    end generate;

    mvb_aligner_g: if META_ALIGN2SOF generate
        mvb_aligner_i : entity work.MVB_ALIGNER
        generic map(
            ITEMS      => REGIONS,
            ITEM_WIDTH => META_WIDTH,
            DEVICE     => DEVICE
        )
        port map(
            CLK        => TX_CLK,
            RESET      => TX_RESET,

            RX_DATA    => slv_array_ser(s_mbuf_mvb_data,REGIONS,META_WIDTH),
            RX_NEW_POS => slv_array_ser(s_mbuf_mvb_new_pos,REGIONS,SOF_INDEX_WIDTH),
            RX_NEW_LIW => s_mbuf_mvb_new_liw,
            RX_FAKE    => s_mbuf_mvb_fake,
            RX_VLD     => s_mbuf_mvb_vld,
            RX_SRC_RDY => s_mbuf_mvb_src_rdy,
            RX_DST_RDY => s_mbuf_mvb_dst_rdy,

            TX_DATA    => TX_MVB_DATA,
            TX_VLD     => TX_MVB_VLD,
            TX_SRC_RDY => TX_MVB_SRC_RDY,
            TX_DST_RDY => TX_MVB_DST_RDY
        );
    else generate
        TX_MVB_DATA        <= slv_array_ser(s_mbuf_mvb_data,REGIONS,META_WIDTH);
        TX_MVB_VLD         <= s_mbuf_mvb_vld;
        TX_MVB_SRC_RDY     <= s_mbuf_mvb_src_rdy;
        s_mbuf_mvb_dst_rdy <= TX_MVB_DST_RDY;
    end generate;

end architecture;
