library IEEE;
use IEEE.std_logic_1164.all;

package dtb_pkg is
    constant DTB_PF0_DATA : std_logic_vector(8*100-1 downto 0) := X"5a590100000000010d994290ab39d6b05c4101005ceb52e300000000d21571da6ddfd6c36acb2615bf684ec2d6d2701fa8b3baea34c962e335a67272f555bed252cd5b0368005d29005b00e0a3e52f74000000160121000236de22690100005a587a37fd";
    constant DTB_VF0_DATA : std_logic_vector(8*100-1 downto 0) := X"5a590100000000010d994290ab39d6b05c4101005ceb52e300000000d21571da6ddfd6c36acb2615bf684ec2d6d2701fa8b3baea34c962e335a67272f555bed252cd5b0368005d29005b00e0a3e52f74000000160121000236de22690100005a587a37fd";
end package dtb_pkg;

package body dtb_pkg is
end dtb_pkg;
