--! testbench.vhd: Testbench of PCIE_MFB2AVST.
--! Copyright (C) 2019 CESNET z. s. p. o.
--! Author(s): Daniel Kondys <xkondy00@vutbr.cz>
--!
--! SPDX-License-Identifier: BSD-3-Clause

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
--! ----------------------------------------------------------------------------
--!                        Entity declaration
--! ----------------------------------------------------------------------------
entity testbench is
end entity testbench;
--! ----------------------------------------------------------------------------
--!                      Architecture declaration
--! ----------------------------------------------------------------------------
architecture behavioral of testbench is
    signal clk            : std_logic;
    signal rst            : std_logic;

    signal mfb_data       : std_logic_vector(511 downto 0);
    signal mfb_meta       : std_logic_vector(15 downto 0);
    signal mfb_sof        : std_logic_vector(1 downto 0);
    signal mfb_eof        : std_logic_vector(1 downto 0);
    signal mfb_eof_pos    : std_logic_vector(5 downto 0);
    signal mfb_src_rdy    : std_logic;
    signal mfb_dst_rdy    : std_logic;

    signal avst_data      : std_logic_vector(511 downto 0);
    signal avst_meta      : std_logic_vector(15 downto 0);
    signal avst_sop       : std_logic_vector(1 downto 0);
    signal avst_eop       : std_logic_vector(1 downto 0);
    signal avst_empty     : std_logic_vector(5 downto 0);
    signal avst_valid     : std_logic_vector(1 downto 0);
    signal avst_dst_rdy   : std_logic;

    constant CLK_PERIOD : time := 10 ns;

    begin
    uut : entity work.PCIE_MFB2AVST
    port map(
        CLK            => clk,
        RST            => rst,

        RX_MFB_DATA    => mfb_data,
        RX_MFB_META    => mfb_meta,
        RX_MFB_SOF     => mfb_sof,
        RX_MFB_EOF     => mfb_eof,
        RX_MFB_EOF_POS => mfb_eof_pos,
        RX_MFB_SRC_RDY => mfb_src_rdy,
        RX_MFB_DST_RDY => mfb_dst_rdy,

        TX_AVST_DATA   => avst_data,
        TX_AVST_META   => avst_meta,
        TX_AVST_SOP    => avst_sop,
        TX_AVST_EOP    => avst_eop,
        TX_AVST_EMPTY  => avst_empty,
        TX_AVST_VALID  => avst_valid,
        TX_AVST_READY  => avst_dst_rdy
    );

    --! generate clk
    clock : process
    begin
       clk <= '1';
       wait for CLK_PERIOD/2;
       clk <= '0';
       wait for CLK_PERIOD/2;
    end process;

    --! generate rst
    reset : process
    begin
       rst <= '1';
       wait for 3*CLK_PERIOD;
       rst <= '0';
       wait;
    end process;

    --! main testbench process for mfb side
    mfb_sim : process
    begin
        mfb_data    <= (others => '0');
        mfb_meta    <= (others => '0');
        mfb_sof     <= (others => '0');
        mfb_eof     <= (others => '0');
        mfb_eof_pos <= (others => '0');
        mfb_src_rdy <= '0';

        wait until rst = '0';

        wait for 0.1*CLK_PERIOD;

     -- =======================================================
     -- testing different SOF and EOF combinations
     -- =======================================================

        mfb_src_rdy <= '1';

        mfb_data <= "00000100000000100110101101010011001001010110101111101100010110000010011100111010000110111010010000001110100100000010011000100010011100110000110000101100011101011110010110100011000101001110111011000100011011111000010111100000110111011100100010110111111101101110100000001111101110000010000100110110010011110001101000111010011110100000001011111100000110111011010111001101100011111110011010100001111111110001100100000100111000100010111001100000111011100100101001100111100010100110001011101101000110110100111111000100";
        mfb_meta <= "0000110100011001";
        mfb_sof <= "11";
        mfb_eof <= "11";
        mfb_eof_pos <= "111110";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if ;

         wait for CLK_PERIOD;

        mfb_data <= "10000010011110110001111101110110110011000010011001001011001110011011011100110000110011110100111100000110100000010110000010001110000001111010011000001101010101011011010100011101010100010011110111000011110100100000001111000100111000100010011001011011010100111001010010001111011000001100000111011000101110110110110010010100111110011111001000111001110111011100011111100000101011010101111001010110001001011110100011000100011101100110010100000011011000100001101110111010101010000011001110011100001100001101111110111111";
        mfb_meta <= "0011010101100000";
        mfb_sof <= "10";
        mfb_eof <= "00";
        mfb_eof_pos <= "000000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if ;

        wait for CLK_PERIOD;

        mfb_data <= "11101100011001000010100011111111111111011100011000110101100000010101101101111100001110111111110010010001101011100101000101011000000110010000010000000100101001110101111101000010001100010110100100000101011101110000100100100111010011110011010001111111010001000111101011110100100100001010001010101101001111000000001010011001100010100011110000111111111010010011110111001010011110110100110011111110000011000010100011100110011111011111110110101100001101011111010011101100000100110000000011100111010000000011101100000011";
        mfb_meta <= "0001100001000110";
        mfb_sof <= "00";
        mfb_eof <= "00";
        mfb_eof_pos <= "000000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "00111100110001000100011000001011000000011010011011011110011011010001101001101000100110001110010101001101110010001001001010001011100001100000000111011001001000001000110101011011111110011110101101011111001011101100100011111001111010001100110111000010000011101111111011100001011101000100001011001100010100101111011100001010001101010000110101001110111000011100000110110101011010010100110111101000110000101110011000001000011100001001111110001101101110110100001000011010001011100010001100111101001010001010111010001111";
        mfb_meta <= "1001101110001011";
        mfb_sof <= "10";
        mfb_eof <= "11";
        mfb_eof_pos <= "010100";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "11010010101100100101010110001010100011001101101010011001111110100110011110100000001111100001110001111100111110001000000000100011100111001010111111100001101010000000010010101000110001000001000101111001000101110111001000111000110010001001100100111101000100011001001001101010110000111111000001011001111011001101010101011010100111011101000000001111001011011100001011011111100011011001000111001110000101101111001100011111110011101110001110111011101010111100000110010100011101101100100011010110111001101110110110010100";
        mfb_meta <= "0001000000100011";
        mfb_sof <= "01";
        mfb_eof <= "10";
        mfb_eof_pos <= "011000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "00010011011100010011001111101101101111111101010101100100111011101001101000101001111100110111000010101101010100000011110001001000110011011000011010101110100110101110111110011001011100100000110100111111000000111101101111011101111101011100011011100010111100100111001111001000110101010110010111000111001100010010011111011111101100000101001100010000100011001101100100111101110100011001111000111111011001101001000001100110011111001001010000010100100101100011011101001000110101101000100101000111011100111001001010000101";
        mfb_meta <= "1111101010001100";
        mfb_sof <= "01";
        mfb_eof <= "00";
        mfb_eof_pos <= "000000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "10100001000010100101000101110010101010011000101000111000001011101000110100110011100100001111000111001001101011010110000000011111001010000100010110000001101100011010111110011111111010111110010110111101110101010010101011011110100011100100000100111110000101110101011011010111010011111111101010111010100111010101101110100101100011101100010110000010011101011110110111110111100000000101010011010100100110111111100111100010101111111111011110010101101000000001110010101110100111011101011010000100101100000001111101001000";
        mfb_meta <= "1001000100111111";
        mfb_sof <= "00";
        mfb_eof <= "10";
        mfb_eof_pos <= "010000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "11011111010111001101010111101100010000001100011000011011011100101001010111011111010000100110101010010001010001110110000000110111110110110010011010111101110001000010110101001100010010111000111001011111111011111010010010111101001101010001011011011001101110010010111100010010100001010101111010101110111111110101100010100111001000000111100110110010010000000101000000101010111101100001000000000011011011100011010110000011111000000100001001010000011110101101100011101010000111100010111110110101111011110100100101100010";
        mfb_meta <= "1001001010001010";
        mfb_sof <= "10";
        mfb_eof <= "10";
        mfb_eof_pos <= "101000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "10110110110110010100010111110110011011111000010010101111011101010001101011010110010100101110001011001101101000110000111101010011001100001110011100001101000101100101100100010000101100100100011100111101000111111101000011011001111010001001011110110001001111110110010110100000010000110110001010011010101011001101000111100110000100101100110111111000001101101010001010101111011110110000000011001000010100101001010101010001111001101101111100001001000011111001101100011010100101101011110101000000110000111010110001010011";
        mfb_meta <= "0101110010101101";
        mfb_sof <= "01";
        mfb_eof <= "01";
        mfb_eof_pos <= "000111";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "00001010000101110101100010001001001001011011001011010011010101011000011111110010000011010000000100010001101000000001011010111011011011100011001101000011111110110010001001100100101111001000101000000000111011101110000010110100100101001000100000100110011000011000110100100010100101001111010100010100110000100000101010101011110111111000010101001000111110001000000101101111010110101010000110100101001100010111110001110110110100111110101111000111001000011111111000101000100101011011001001010000011001011111101110110001";
        mfb_meta <= "1100110011001001";
        mfb_sof <= "10";
        mfb_eof <= "00";
        mfb_eof_pos <= "000000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "10110011010001010101010011100111010110000110010011111101001010010010000100010101000000110101010011000101101100010110100011001100101100101100100001110010101110110101100001001000010011011010111100101100010000100101110110011100010100110001010000100101100100110100100111111001110111101001110111111000010010101010010011010110010011011010001100010011011101111001111010110101101000011101111111001100000100010000110011111111000100000111010110110101100111110110001110011111001110100000110010110101001101100110001110011010";
        mfb_meta <= "1010011011000011";
        mfb_sof <= "10";
        mfb_eof <= "01";
        mfb_eof_pos <= "000101";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "10011100000011011001000111010111101010001011001010000110011110001001011011101011011100011000010011001011011100010001000010110011110101010100010100010001011110110001000000111101101111011010010101111110011000000111011110011110001000000110011001000111000111001110000101001011010100011011001010000001111010110111100100111110100001011111101110111010101110011101001011001000110001011101100100100011010110101000111101111101100010010001111001101100100110100000111101011001100111101110111100010011010100001010111010111111";
        mfb_meta <= "1100000100111111";
        mfb_sof <= "00";
        mfb_eof <= "01";
        mfb_eof_pos <= "000111";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        -- =======================================================
        -- testing different src_rdy and dst_rdy combinations
        -- =======================================================

        mfb_src_rdy <= '1'; -- this is already set, just a reminder
        -- avst_dst_rdy <= '0'; -- this is set in the next process, just as a clarification

        mfb_data <= "10100101001000111100100110111100010111110111000111100000101011001011101110010001010100000010000001110110111100000001100001110101000111100010100101111010001010110000000010000010101100011110000100110101100110100100000000001000001110111010110101000110101111011101000011110111111101010011000001110111110101100101111101110010000110111101000111010101010110000011001001100000111011000100000100100010101000110110101000111101000101011111100110110011111110010000001001110001010011111011011110101001110110110001011010101111";
        mfb_meta <= "1101100100000010";
        mfb_sof <= "11";
        mfb_eof <= "11";
        mfb_eof_pos <= "011111";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "10100111011100000011011110010110011011011101101111110010011111101011110011110001100011000000011100101000010101010101010111011011110010011100111011000110111110001010000001011101001010111010010100110000000101011110010110101110000010010111010001111000001111000011001101010000110011100001100011111001001111011101110101000101110101100110011001101101010110000110010010100000010101001000001100100010100110111000111000000110101010001001011010100010110101101011100101111011001000011001101110101011011011000111111111010010";
        mfb_meta <= "1110111100000000";
        mfb_sof <= "11";
        mfb_eof <= "11";
        mfb_eof_pos <= "011111";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "11101100011001000010100011111111100111011100011000110101100000010101101101111100001110111111110010010001101011100101000101011000000110010000010000000100101001110101111101000010001100010110100100000101011101110000100100100111010011110011010001111111010001000111101011110100100100001010001010101101001111000000001010011001100010100011110000111111111010010011110111001010011110110100110011111110000011000010100011100110011111011111110110101100001101011111010011101100000100110000000011100111010000000011101100000011";
        mfb_meta <= "1011101011111111";
        mfb_sof <= "01";
        mfb_eof <= "10";
        mfb_eof_pos <= "101000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_src_rdy <= '1';

        mfb_data <= "10101010100000011001110000000011101100011110011010010101110011101100001110110110101100100111001010001111000111111110000101110010101000011000110110000100001111111111010111001011001011100101010011100111000101010011000011101101100110001101111100011011111100110011010111000000101011100100011010101111101011100100000010101010100010111011110111111101000100110010011101000000110011000101011101011111110011111100111001111110110010101110100111100010100101111001100111100100011101010001010110110100000111011000110101011010";
        mfb_meta <= "0111000010011110";
        mfb_sof <= "01";
        mfb_eof <= "10";
        mfb_eof_pos <= "010000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_data <= "00101011100011001010100011010110000001001010111101011101100101110101100011111001000010010000011111111100100110101101100010101010111001011011000011001101100001010110001111100101000001011100010010111100011010110110010100010011111101100100011010001011001010001100100110001110110111001011110010100000111110010110111001010000001011000100001110000010101110110001010011011000010010100000010110010101101011011010010100010000000000010111111010010011001111111000001100100000001000100000101010010101111011010101100100010010";
        mfb_meta <= "1011100000000011";
        mfb_sof <= "01";
        mfb_eof <= "10";
        mfb_eof_pos <= "110000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_src_rdy <= '0';

        mfb_data <= "11001111101111110011011010001011110111000110011011100111011110010000011110010110010101100011100110010100000101111111111110110011100101111010000001110111110101011101110101111110011111100110011000110000101000010001101111011101011010011110010101100110000110010011011010000001111101010001100100100111010101000001101011111010010100000101111111001110001111100000000100001111011110101000011010010011101101001011100101111001101000011110111100111110010001010110000111100001010001010000000010011100101111101101011001110100";
        mfb_meta <= "0010101001110111";
        mfb_sof <= "01";
        mfb_eof <= "10";
        mfb_eof_pos <= "011000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_src_rdy <= '0';

        mfb_data <= "01010011011001111010010111010101101100110100001010110001001010100111010001111001111010011010100011100001110100111001111010100101101010110101010100001001111111100011100000011110111010100000111000010010011010111001100111100100001000011110110011101110000101010001011100100111010110111001010001010011100010100100111001011111011000011111001011100011111011011101111111000011001010110000110111010101101001000111011101000001001010110110010110110111011010101001010001010010001001011011111010111010111111100010011011001011";
        mfb_meta <= "1100101001010100";
        mfb_sof <= "01";
        mfb_eof <= "10";
        mfb_eof_pos <= "001000";
        if mfb_dst_rdy = '0' then
            wait until mfb_dst_rdy = '1';
            wait for 0.1*CLK_PERIOD;
        end if;

        wait for CLK_PERIOD;

        mfb_src_rdy <= '1';

        wait;
    end process;

    --! main testbench process for avst side
    avst_sim : process
    begin
        avst_dst_rdy <= '0';

        wait until rst = '0';

        wait for 0.1*CLK_PERIOD;

        avst_dst_rdy <= '1';

        wait for 13*CLK_PERIOD;

        avst_dst_rdy <= '0';

        wait for 4*CLK_PERIOD;

        avst_dst_rdy <= '1';

        wait for 3*CLK_PERIOD;

        avst_dst_rdy <= '0';

        wait for CLK_PERIOD;

        avst_dst_rdy <= '1';

        wait;
    end process;

end architecture behavioral;